module PixelOffreg( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [31:0] io_start_x, // @[:@6.4]
  input  [31:0] io_start_y, // @[:@6.4]
  input  [31:0] io_del_x, // @[:@6.4]
  input  [31:0] io_del_y, // @[:@6.4]
  output [31:0] io_offset_x_0, // @[:@6.4]
  output [31:0] io_offset_x_1, // @[:@6.4]
  output [31:0] io_offset_x_2, // @[:@6.4]
  output [31:0] io_offset_x_3, // @[:@6.4]
  output [31:0] io_offset_x_4, // @[:@6.4]
  output [31:0] io_offset_x_5, // @[:@6.4]
  output [31:0] io_offset_x_6, // @[:@6.4]
  output [31:0] io_offset_x_7, // @[:@6.4]
  output [31:0] io_offset_x_8, // @[:@6.4]
  output [31:0] io_offset_x_9, // @[:@6.4]
  output [31:0] io_offset_x_10, // @[:@6.4]
  output [31:0] io_offset_x_11, // @[:@6.4]
  output [31:0] io_offset_x_12, // @[:@6.4]
  output [31:0] io_offset_x_13, // @[:@6.4]
  output [31:0] io_offset_x_14, // @[:@6.4]
  output [31:0] io_offset_x_15, // @[:@6.4]
  output [31:0] io_offset_y_0, // @[:@6.4]
  output [31:0] io_offset_y_1, // @[:@6.4]
  output [31:0] io_offset_y_2, // @[:@6.4]
  output [31:0] io_offset_y_3, // @[:@6.4]
  output [31:0] io_offset_y_4, // @[:@6.4]
  output [31:0] io_offset_y_5, // @[:@6.4]
  output [31:0] io_offset_y_6, // @[:@6.4]
  output [31:0] io_offset_y_7, // @[:@6.4]
  output [31:0] io_offset_y_8, // @[:@6.4]
  output [31:0] io_offset_y_9, // @[:@6.4]
  output [31:0] io_offset_y_10, // @[:@6.4]
  output [31:0] io_offset_y_11, // @[:@6.4]
  output [31:0] io_offset_y_12, // @[:@6.4]
  output [31:0] io_offset_y_13, // @[:@6.4]
  output [31:0] io_offset_y_14, // @[:@6.4]
  output [31:0] io_offset_y_15, // @[:@6.4]
  output [31:0] io_vld // @[:@6.4]
);
  wire [31:0] _T_99; // @[offreg.scala 18:50:@8.4]
  wire [31:0] _T_100; // @[offreg.scala 18:82:@9.4]
  wire [31:0] _T_101; // @[offreg.scala 19:46:@10.4]
  wire [31:0] _T_102; // @[offreg.scala 19:76:@11.4]
  wire [31:0] _T_103; // @[offreg.scala 65:23:@12.4]
  wire [27:0] _T_104; // @[offreg.scala 65:26:@13.4]
  wire [28:0] _T_105; // @[offreg.scala 65:32:@14.4]
  wire [28:0] _T_106; // @[offreg.scala 65:52:@15.4]
  wire [22:0] _T_107; // @[offreg.scala 65:60:@16.4]
  wire [31:0] _T_108; // @[offreg.scala 66:23:@17.4]
  wire [27:0] _T_109; // @[offreg.scala 66:26:@18.4]
  wire [28:0] _T_110; // @[offreg.scala 66:32:@19.4]
  wire [28:0] _T_111; // @[offreg.scala 66:52:@20.4]
  wire [22:0] _T_112; // @[offreg.scala 66:60:@21.4]
  wire [31:0] _GEN_0; // @[offreg.scala 59:15:@22.4]
  wire [32:0] _T_113; // @[offreg.scala 59:15:@22.4]
  wire [31:0] _T_114; // @[offreg.scala 59:15:@23.4]
  wire [31:0] _T_115; // @[offreg.scala 59:15:@24.4]
  wire [31:0] _GEN_1; // @[offreg.scala 60:15:@25.4]
  wire [32:0] _T_116; // @[offreg.scala 60:15:@25.4]
  wire [31:0] _T_117; // @[offreg.scala 60:15:@26.4]
  wire [31:0] _T_118; // @[offreg.scala 60:15:@27.4]
  wire [29:0] _T_121; // @[offreg.scala 65:32:@30.4]
  wire [29:0] _T_122; // @[offreg.scala 65:52:@31.4]
  wire [23:0] _T_123; // @[offreg.scala 65:60:@32.4]
  wire [29:0] _T_126; // @[offreg.scala 66:32:@35.4]
  wire [29:0] _T_127; // @[offreg.scala 66:52:@36.4]
  wire [23:0] _T_128; // @[offreg.scala 66:60:@37.4]
  wire [31:0] _GEN_2; // @[offreg.scala 59:15:@38.4]
  wire [32:0] _T_129; // @[offreg.scala 59:15:@38.4]
  wire [31:0] _T_130; // @[offreg.scala 59:15:@39.4]
  wire [31:0] _T_131; // @[offreg.scala 59:15:@40.4]
  wire [31:0] _GEN_3; // @[offreg.scala 60:15:@41.4]
  wire [32:0] _T_132; // @[offreg.scala 60:15:@41.4]
  wire [31:0] _T_133; // @[offreg.scala 60:15:@42.4]
  wire [31:0] _T_134; // @[offreg.scala 60:15:@43.4]
  wire [30:0] _T_137; // @[offreg.scala 65:32:@46.4]
  wire [30:0] _T_138; // @[offreg.scala 65:52:@47.4]
  wire [24:0] _T_139; // @[offreg.scala 65:60:@48.4]
  wire [30:0] _T_142; // @[offreg.scala 66:32:@51.4]
  wire [30:0] _T_143; // @[offreg.scala 66:52:@52.4]
  wire [24:0] _T_144; // @[offreg.scala 66:60:@53.4]
  wire [31:0] _GEN_4; // @[offreg.scala 59:15:@54.4]
  wire [32:0] _T_145; // @[offreg.scala 59:15:@54.4]
  wire [31:0] _T_146; // @[offreg.scala 59:15:@55.4]
  wire [31:0] _T_147; // @[offreg.scala 59:15:@56.4]
  wire [31:0] _GEN_5; // @[offreg.scala 60:15:@57.4]
  wire [32:0] _T_148; // @[offreg.scala 60:15:@57.4]
  wire [31:0] _T_149; // @[offreg.scala 60:15:@58.4]
  wire [31:0] _T_150; // @[offreg.scala 60:15:@59.4]
  wire [30:0] _T_153; // @[offreg.scala 65:32:@62.4]
  wire [30:0] _T_154; // @[offreg.scala 65:52:@63.4]
  wire [24:0] _T_155; // @[offreg.scala 65:60:@64.4]
  wire [30:0] _T_158; // @[offreg.scala 66:32:@67.4]
  wire [30:0] _T_159; // @[offreg.scala 66:52:@68.4]
  wire [24:0] _T_160; // @[offreg.scala 66:60:@69.4]
  wire [31:0] _GEN_6; // @[offreg.scala 59:15:@70.4]
  wire [32:0] _T_161; // @[offreg.scala 59:15:@70.4]
  wire [31:0] _T_162; // @[offreg.scala 59:15:@71.4]
  wire [31:0] _T_163; // @[offreg.scala 59:15:@72.4]
  wire [31:0] _GEN_7; // @[offreg.scala 60:15:@73.4]
  wire [32:0] _T_164; // @[offreg.scala 60:15:@73.4]
  wire [31:0] _T_165; // @[offreg.scala 60:15:@74.4]
  wire [31:0] _T_166; // @[offreg.scala 60:15:@75.4]
  wire [31:0] _T_169; // @[offreg.scala 65:32:@78.4]
  wire [31:0] _T_170; // @[offreg.scala 65:52:@79.4]
  wire [25:0] _T_171; // @[offreg.scala 65:60:@80.4]
  wire [31:0] _T_174; // @[offreg.scala 66:32:@83.4]
  wire [31:0] _T_175; // @[offreg.scala 66:52:@84.4]
  wire [25:0] _T_176; // @[offreg.scala 66:60:@85.4]
  wire [31:0] _GEN_8; // @[offreg.scala 59:15:@86.4]
  wire [32:0] _T_177; // @[offreg.scala 59:15:@86.4]
  wire [31:0] _T_178; // @[offreg.scala 59:15:@87.4]
  wire [31:0] _T_179; // @[offreg.scala 59:15:@88.4]
  wire [31:0] _GEN_9; // @[offreg.scala 60:15:@89.4]
  wire [32:0] _T_180; // @[offreg.scala 60:15:@89.4]
  wire [31:0] _T_181; // @[offreg.scala 60:15:@90.4]
  wire [31:0] _T_182; // @[offreg.scala 60:15:@91.4]
  wire [31:0] _T_185; // @[offreg.scala 65:32:@94.4]
  wire [31:0] _T_186; // @[offreg.scala 65:52:@95.4]
  wire [25:0] _T_187; // @[offreg.scala 65:60:@96.4]
  wire [31:0] _T_190; // @[offreg.scala 66:32:@99.4]
  wire [31:0] _T_191; // @[offreg.scala 66:52:@100.4]
  wire [25:0] _T_192; // @[offreg.scala 66:60:@101.4]
  wire [31:0] _GEN_10; // @[offreg.scala 59:15:@102.4]
  wire [32:0] _T_193; // @[offreg.scala 59:15:@102.4]
  wire [31:0] _T_194; // @[offreg.scala 59:15:@103.4]
  wire [31:0] _T_195; // @[offreg.scala 59:15:@104.4]
  wire [31:0] _GEN_11; // @[offreg.scala 60:15:@105.4]
  wire [32:0] _T_196; // @[offreg.scala 60:15:@105.4]
  wire [31:0] _T_197; // @[offreg.scala 60:15:@106.4]
  wire [31:0] _T_198; // @[offreg.scala 60:15:@107.4]
  wire [31:0] _T_201; // @[offreg.scala 65:32:@110.4]
  wire [31:0] _T_202; // @[offreg.scala 65:52:@111.4]
  wire [25:0] _T_203; // @[offreg.scala 65:60:@112.4]
  wire [31:0] _T_206; // @[offreg.scala 66:32:@115.4]
  wire [31:0] _T_207; // @[offreg.scala 66:52:@116.4]
  wire [25:0] _T_208; // @[offreg.scala 66:60:@117.4]
  wire [31:0] _GEN_12; // @[offreg.scala 59:15:@118.4]
  wire [32:0] _T_209; // @[offreg.scala 59:15:@118.4]
  wire [31:0] _T_210; // @[offreg.scala 59:15:@119.4]
  wire [31:0] _T_211; // @[offreg.scala 59:15:@120.4]
  wire [31:0] _GEN_13; // @[offreg.scala 60:15:@121.4]
  wire [32:0] _T_212; // @[offreg.scala 60:15:@121.4]
  wire [31:0] _T_213; // @[offreg.scala 60:15:@122.4]
  wire [31:0] _T_214; // @[offreg.scala 60:15:@123.4]
  wire [31:0] _T_217; // @[offreg.scala 65:32:@126.4]
  wire [31:0] _T_218; // @[offreg.scala 65:52:@127.4]
  wire [25:0] _T_219; // @[offreg.scala 65:60:@128.4]
  wire [31:0] _T_222; // @[offreg.scala 66:32:@131.4]
  wire [31:0] _T_223; // @[offreg.scala 66:52:@132.4]
  wire [25:0] _T_224; // @[offreg.scala 66:60:@133.4]
  wire [31:0] _GEN_14; // @[offreg.scala 59:15:@134.4]
  wire [32:0] _T_225; // @[offreg.scala 59:15:@134.4]
  wire [31:0] _T_226; // @[offreg.scala 59:15:@135.4]
  wire [31:0] _T_227; // @[offreg.scala 59:15:@136.4]
  wire [31:0] _GEN_15; // @[offreg.scala 60:15:@137.4]
  wire [32:0] _T_228; // @[offreg.scala 60:15:@137.4]
  wire [31:0] _T_229; // @[offreg.scala 60:15:@138.4]
  wire [31:0] _T_230; // @[offreg.scala 60:15:@139.4]
  wire [32:0] _T_233; // @[offreg.scala 65:32:@142.4]
  wire [32:0] _T_234; // @[offreg.scala 65:52:@143.4]
  wire [26:0] _T_235; // @[offreg.scala 65:60:@144.4]
  wire [32:0] _T_238; // @[offreg.scala 66:32:@147.4]
  wire [32:0] _T_239; // @[offreg.scala 66:52:@148.4]
  wire [26:0] _T_240; // @[offreg.scala 66:60:@149.4]
  wire [31:0] _GEN_16; // @[offreg.scala 59:15:@150.4]
  wire [32:0] _T_241; // @[offreg.scala 59:15:@150.4]
  wire [31:0] _T_242; // @[offreg.scala 59:15:@151.4]
  wire [31:0] _T_243; // @[offreg.scala 59:15:@152.4]
  wire [31:0] _GEN_17; // @[offreg.scala 60:15:@153.4]
  wire [32:0] _T_244; // @[offreg.scala 60:15:@153.4]
  wire [31:0] _T_245; // @[offreg.scala 60:15:@154.4]
  wire [31:0] _T_246; // @[offreg.scala 60:15:@155.4]
  wire [32:0] _T_249; // @[offreg.scala 65:32:@158.4]
  wire [32:0] _T_250; // @[offreg.scala 65:52:@159.4]
  wire [26:0] _T_251; // @[offreg.scala 65:60:@160.4]
  wire [32:0] _T_254; // @[offreg.scala 66:32:@163.4]
  wire [32:0] _T_255; // @[offreg.scala 66:52:@164.4]
  wire [26:0] _T_256; // @[offreg.scala 66:60:@165.4]
  wire [31:0] _GEN_18; // @[offreg.scala 59:15:@166.4]
  wire [32:0] _T_257; // @[offreg.scala 59:15:@166.4]
  wire [31:0] _T_258; // @[offreg.scala 59:15:@167.4]
  wire [31:0] _T_259; // @[offreg.scala 59:15:@168.4]
  wire [31:0] _GEN_19; // @[offreg.scala 60:15:@169.4]
  wire [32:0] _T_260; // @[offreg.scala 60:15:@169.4]
  wire [31:0] _T_261; // @[offreg.scala 60:15:@170.4]
  wire [31:0] _T_262; // @[offreg.scala 60:15:@171.4]
  wire [32:0] _T_265; // @[offreg.scala 65:32:@174.4]
  wire [32:0] _T_266; // @[offreg.scala 65:52:@175.4]
  wire [26:0] _T_267; // @[offreg.scala 65:60:@176.4]
  wire [32:0] _T_270; // @[offreg.scala 66:32:@179.4]
  wire [32:0] _T_271; // @[offreg.scala 66:52:@180.4]
  wire [26:0] _T_272; // @[offreg.scala 66:60:@181.4]
  wire [31:0] _GEN_20; // @[offreg.scala 59:15:@182.4]
  wire [32:0] _T_273; // @[offreg.scala 59:15:@182.4]
  wire [31:0] _T_274; // @[offreg.scala 59:15:@183.4]
  wire [31:0] _T_275; // @[offreg.scala 59:15:@184.4]
  wire [31:0] _GEN_21; // @[offreg.scala 60:15:@185.4]
  wire [32:0] _T_276; // @[offreg.scala 60:15:@185.4]
  wire [31:0] _T_277; // @[offreg.scala 60:15:@186.4]
  wire [31:0] _T_278; // @[offreg.scala 60:15:@187.4]
  wire [32:0] _T_281; // @[offreg.scala 65:32:@190.4]
  wire [32:0] _T_282; // @[offreg.scala 65:52:@191.4]
  wire [26:0] _T_283; // @[offreg.scala 65:60:@192.4]
  wire [32:0] _T_286; // @[offreg.scala 66:32:@195.4]
  wire [32:0] _T_287; // @[offreg.scala 66:52:@196.4]
  wire [26:0] _T_288; // @[offreg.scala 66:60:@197.4]
  wire [31:0] _GEN_22; // @[offreg.scala 59:15:@198.4]
  wire [32:0] _T_289; // @[offreg.scala 59:15:@198.4]
  wire [31:0] _T_290; // @[offreg.scala 59:15:@199.4]
  wire [31:0] _T_291; // @[offreg.scala 59:15:@200.4]
  wire [31:0] _GEN_23; // @[offreg.scala 60:15:@201.4]
  wire [32:0] _T_292; // @[offreg.scala 60:15:@201.4]
  wire [31:0] _T_293; // @[offreg.scala 60:15:@202.4]
  wire [31:0] _T_294; // @[offreg.scala 60:15:@203.4]
  wire [32:0] _T_297; // @[offreg.scala 65:32:@206.4]
  wire [32:0] _T_298; // @[offreg.scala 65:52:@207.4]
  wire [26:0] _T_299; // @[offreg.scala 65:60:@208.4]
  wire [32:0] _T_302; // @[offreg.scala 66:32:@211.4]
  wire [32:0] _T_303; // @[offreg.scala 66:52:@212.4]
  wire [26:0] _T_304; // @[offreg.scala 66:60:@213.4]
  wire [31:0] _GEN_24; // @[offreg.scala 59:15:@214.4]
  wire [32:0] _T_305; // @[offreg.scala 59:15:@214.4]
  wire [31:0] _T_306; // @[offreg.scala 59:15:@215.4]
  wire [31:0] _T_307; // @[offreg.scala 59:15:@216.4]
  wire [31:0] _GEN_25; // @[offreg.scala 60:15:@217.4]
  wire [32:0] _T_308; // @[offreg.scala 60:15:@217.4]
  wire [31:0] _T_309; // @[offreg.scala 60:15:@218.4]
  wire [31:0] _T_310; // @[offreg.scala 60:15:@219.4]
  wire [32:0] _T_313; // @[offreg.scala 65:32:@222.4]
  wire [32:0] _T_314; // @[offreg.scala 65:52:@223.4]
  wire [26:0] _T_315; // @[offreg.scala 65:60:@224.4]
  wire [32:0] _T_318; // @[offreg.scala 66:32:@227.4]
  wire [32:0] _T_319; // @[offreg.scala 66:52:@228.4]
  wire [26:0] _T_320; // @[offreg.scala 66:60:@229.4]
  wire [31:0] _GEN_26; // @[offreg.scala 59:15:@230.4]
  wire [32:0] _T_321; // @[offreg.scala 59:15:@230.4]
  wire [31:0] _T_322; // @[offreg.scala 59:15:@231.4]
  wire [31:0] _T_323; // @[offreg.scala 59:15:@232.4]
  wire [31:0] _GEN_27; // @[offreg.scala 60:15:@233.4]
  wire [32:0] _T_324; // @[offreg.scala 60:15:@233.4]
  wire [31:0] _T_325; // @[offreg.scala 60:15:@234.4]
  wire [31:0] _T_326; // @[offreg.scala 60:15:@235.4]
  wire [32:0] _T_329; // @[offreg.scala 65:32:@238.4]
  wire [32:0] _T_330; // @[offreg.scala 65:52:@239.4]
  wire [26:0] _T_331; // @[offreg.scala 65:60:@240.4]
  wire [32:0] _T_334; // @[offreg.scala 66:32:@243.4]
  wire [32:0] _T_335; // @[offreg.scala 66:52:@244.4]
  wire [26:0] _T_336; // @[offreg.scala 66:60:@245.4]
  wire [31:0] _GEN_28; // @[offreg.scala 59:15:@246.4]
  wire [32:0] _T_337; // @[offreg.scala 59:15:@246.4]
  wire [31:0] _T_338; // @[offreg.scala 59:15:@247.4]
  wire [31:0] _T_339; // @[offreg.scala 59:15:@248.4]
  wire [31:0] _GEN_29; // @[offreg.scala 60:15:@249.4]
  wire [32:0] _T_340; // @[offreg.scala 60:15:@249.4]
  wire [31:0] _T_341; // @[offreg.scala 60:15:@250.4]
  wire [31:0] _T_342; // @[offreg.scala 60:15:@251.4]
  wire [32:0] _T_345; // @[offreg.scala 65:32:@254.4]
  wire [32:0] _T_346; // @[offreg.scala 65:52:@255.4]
  wire [26:0] _T_347; // @[offreg.scala 65:60:@256.4]
  wire [32:0] _T_350; // @[offreg.scala 66:32:@259.4]
  wire [32:0] _T_351; // @[offreg.scala 66:52:@260.4]
  wire [26:0] _T_352; // @[offreg.scala 66:60:@261.4]
  wire [31:0] _GEN_30; // @[offreg.scala 59:15:@262.4]
  wire [32:0] _T_353; // @[offreg.scala 59:15:@262.4]
  wire [31:0] _T_354; // @[offreg.scala 59:15:@263.4]
  wire [31:0] _T_355; // @[offreg.scala 59:15:@264.4]
  wire [31:0] _GEN_31; // @[offreg.scala 60:15:@265.4]
  wire [32:0] _T_356; // @[offreg.scala 60:15:@265.4]
  wire [31:0] _T_357; // @[offreg.scala 60:15:@266.4]
  wire [31:0] _T_358; // @[offreg.scala 60:15:@267.4]
  wire [32:0] _T_393; // @[offreg.scala 59:15:@332.4]
  wire [31:0] _T_394; // @[offreg.scala 59:15:@333.4]
  wire [31:0] _T_395; // @[offreg.scala 59:15:@334.4]
  wire [32:0] _T_396; // @[offreg.scala 60:15:@335.4]
  wire [31:0] _T_397; // @[offreg.scala 60:15:@336.4]
  wire [31:0] _T_398; // @[offreg.scala 60:15:@337.4]
  wire  _T_399; // @[offreg.scala 70:12:@338.4]
  wire  _T_400; // @[offreg.scala 70:26:@339.4]
  wire  vld_0; // @[offreg.scala 70:20:@340.4]
  wire  _T_401; // @[offreg.scala 70:12:@341.4]
  wire  _T_402; // @[offreg.scala 70:26:@342.4]
  wire  vld_1; // @[offreg.scala 70:20:@343.4]
  wire  _T_403; // @[offreg.scala 70:12:@344.4]
  wire  _T_404; // @[offreg.scala 70:26:@345.4]
  wire  vld_2; // @[offreg.scala 70:20:@346.4]
  wire  _T_405; // @[offreg.scala 70:12:@347.4]
  wire  _T_406; // @[offreg.scala 70:26:@348.4]
  wire  vld_3; // @[offreg.scala 70:20:@349.4]
  wire  _T_407; // @[offreg.scala 70:12:@350.4]
  wire  _T_408; // @[offreg.scala 70:26:@351.4]
  wire  vld_4; // @[offreg.scala 70:20:@352.4]
  wire  _T_409; // @[offreg.scala 70:12:@353.4]
  wire  _T_410; // @[offreg.scala 70:26:@354.4]
  wire  vld_5; // @[offreg.scala 70:20:@355.4]
  wire  _T_411; // @[offreg.scala 70:12:@356.4]
  wire  _T_412; // @[offreg.scala 70:26:@357.4]
  wire  vld_6; // @[offreg.scala 70:20:@358.4]
  wire  _T_413; // @[offreg.scala 70:12:@359.4]
  wire  _T_414; // @[offreg.scala 70:26:@360.4]
  wire  vld_7; // @[offreg.scala 70:20:@361.4]
  wire  _T_415; // @[offreg.scala 70:12:@362.4]
  wire  _T_416; // @[offreg.scala 70:26:@363.4]
  wire  vld_8; // @[offreg.scala 70:20:@364.4]
  wire  _T_417; // @[offreg.scala 70:12:@365.4]
  wire  _T_418; // @[offreg.scala 70:26:@366.4]
  wire  vld_9; // @[offreg.scala 70:20:@367.4]
  wire  _T_419; // @[offreg.scala 70:12:@368.4]
  wire  _T_420; // @[offreg.scala 70:26:@369.4]
  wire  vld_10; // @[offreg.scala 70:20:@370.4]
  wire  _T_421; // @[offreg.scala 70:12:@371.4]
  wire  _T_422; // @[offreg.scala 70:26:@372.4]
  wire  vld_11; // @[offreg.scala 70:20:@373.4]
  wire  _T_423; // @[offreg.scala 70:12:@374.4]
  wire  _T_424; // @[offreg.scala 70:26:@375.4]
  wire  vld_12; // @[offreg.scala 70:20:@376.4]
  wire  _T_425; // @[offreg.scala 70:12:@377.4]
  wire  _T_426; // @[offreg.scala 70:26:@378.4]
  wire  vld_13; // @[offreg.scala 70:20:@379.4]
  wire  _T_427; // @[offreg.scala 70:12:@380.4]
  wire  _T_428; // @[offreg.scala 70:26:@381.4]
  wire  vld_14; // @[offreg.scala 70:20:@382.4]
  wire  _T_429; // @[offreg.scala 70:12:@383.4]
  wire  _T_430; // @[offreg.scala 70:26:@384.4]
  wire  vld_15; // @[offreg.scala 70:20:@385.4]
  wire [1:0] _GEN_32; // @[offreg.scala 32:52:@387.4]
  wire [1:0] _T_432; // @[offreg.scala 32:52:@387.4]
  wire [2:0] _GEN_33; // @[offreg.scala 32:52:@388.4]
  wire [2:0] _T_433; // @[offreg.scala 32:52:@388.4]
  wire [3:0] _GEN_34; // @[offreg.scala 32:52:@389.4]
  wire [3:0] _T_434; // @[offreg.scala 32:52:@389.4]
  wire [4:0] _GEN_35; // @[offreg.scala 32:52:@390.4]
  wire [4:0] _T_435; // @[offreg.scala 32:52:@390.4]
  wire [5:0] _GEN_36; // @[offreg.scala 32:52:@391.4]
  wire [5:0] _T_436; // @[offreg.scala 32:52:@391.4]
  wire [6:0] _GEN_37; // @[offreg.scala 32:52:@392.4]
  wire [6:0] _T_437; // @[offreg.scala 32:52:@392.4]
  wire [7:0] _GEN_38; // @[offreg.scala 32:52:@393.4]
  wire [7:0] _T_438; // @[offreg.scala 32:52:@393.4]
  wire [8:0] _GEN_39; // @[offreg.scala 32:52:@394.4]
  wire [8:0] _T_439; // @[offreg.scala 32:52:@394.4]
  wire [9:0] _GEN_40; // @[offreg.scala 32:52:@395.4]
  wire [9:0] _T_440; // @[offreg.scala 32:52:@395.4]
  wire [10:0] _GEN_41; // @[offreg.scala 32:52:@396.4]
  wire [10:0] _T_441; // @[offreg.scala 32:52:@396.4]
  wire [11:0] _GEN_42; // @[offreg.scala 32:52:@397.4]
  wire [11:0] _T_442; // @[offreg.scala 32:52:@397.4]
  wire [12:0] _GEN_43; // @[offreg.scala 32:52:@398.4]
  wire [12:0] _T_443; // @[offreg.scala 32:52:@398.4]
  wire [13:0] _GEN_44; // @[offreg.scala 32:52:@399.4]
  wire [13:0] _T_444; // @[offreg.scala 32:52:@399.4]
  wire [14:0] _GEN_45; // @[offreg.scala 32:52:@400.4]
  wire [14:0] _T_445; // @[offreg.scala 32:52:@400.4]
  wire [15:0] _GEN_46; // @[offreg.scala 32:52:@401.4]
  wire [15:0] _T_446; // @[offreg.scala 32:52:@401.4]
  wire [1:0] _GEN_47; // @[offreg.scala 32:74:@403.4]
  wire [1:0] _T_449; // @[offreg.scala 32:74:@403.4]
  wire [2:0] _GEN_48; // @[offreg.scala 32:74:@404.4]
  wire [2:0] _T_450; // @[offreg.scala 32:74:@404.4]
  wire [3:0] _GEN_49; // @[offreg.scala 32:74:@405.4]
  wire [3:0] _T_451; // @[offreg.scala 32:74:@405.4]
  wire [4:0] _GEN_50; // @[offreg.scala 32:74:@406.4]
  wire [4:0] _T_452; // @[offreg.scala 32:74:@406.4]
  wire [5:0] _GEN_51; // @[offreg.scala 32:74:@407.4]
  wire [5:0] _T_453; // @[offreg.scala 32:74:@407.4]
  wire [6:0] _GEN_52; // @[offreg.scala 32:74:@408.4]
  wire [6:0] _T_454; // @[offreg.scala 32:74:@408.4]
  wire [7:0] _GEN_53; // @[offreg.scala 32:74:@409.4]
  wire [7:0] _T_455; // @[offreg.scala 32:74:@409.4]
  wire [8:0] _GEN_54; // @[offreg.scala 32:74:@410.4]
  wire [8:0] _T_456; // @[offreg.scala 32:74:@410.4]
  wire [9:0] _GEN_55; // @[offreg.scala 32:74:@411.4]
  wire [9:0] _T_457; // @[offreg.scala 32:74:@411.4]
  wire [10:0] _GEN_56; // @[offreg.scala 32:74:@412.4]
  wire [10:0] _T_458; // @[offreg.scala 32:74:@412.4]
  wire [11:0] _GEN_57; // @[offreg.scala 32:74:@413.4]
  wire [11:0] _T_459; // @[offreg.scala 32:74:@413.4]
  wire [12:0] _GEN_58; // @[offreg.scala 32:74:@414.4]
  wire [12:0] _T_460; // @[offreg.scala 32:74:@414.4]
  wire [13:0] _GEN_59; // @[offreg.scala 32:74:@415.4]
  wire [13:0] _T_461; // @[offreg.scala 32:74:@415.4]
  wire [14:0] _GEN_60; // @[offreg.scala 32:74:@416.4]
  wire [14:0] _T_462; // @[offreg.scala 32:74:@416.4]
  wire [15:0] _GEN_61; // @[offreg.scala 32:74:@417.4]
  wire [15:0] _T_463; // @[offreg.scala 32:74:@417.4]
  assign _T_99 = $signed(io_start_x); // @[offreg.scala 18:50:@8.4]
  assign _T_100 = $signed(io_start_y); // @[offreg.scala 18:82:@9.4]
  assign _T_101 = $signed(io_del_x); // @[offreg.scala 19:46:@10.4]
  assign _T_102 = $signed(io_del_y); // @[offreg.scala 19:76:@11.4]
  assign _T_103 = $signed(_T_101); // @[offreg.scala 65:23:@12.4]
  assign _T_104 = _T_103[31:4]; // @[offreg.scala 65:26:@13.4]
  assign _T_105 = $signed(_T_104) * $signed(28'sh0); // @[offreg.scala 65:32:@14.4]
  assign _T_106 = $signed(_T_105); // @[offreg.scala 65:52:@15.4]
  assign _T_107 = _T_106[28:6]; // @[offreg.scala 65:60:@16.4]
  assign _T_108 = $signed(_T_102); // @[offreg.scala 66:23:@17.4]
  assign _T_109 = _T_108[31:4]; // @[offreg.scala 66:26:@18.4]
  assign _T_110 = $signed(_T_109) * $signed(28'sh0); // @[offreg.scala 66:32:@19.4]
  assign _T_111 = $signed(_T_110); // @[offreg.scala 66:52:@20.4]
  assign _T_112 = _T_111[28:6]; // @[offreg.scala 66:60:@21.4]
  assign _GEN_0 = {{9{_T_107[22]}},_T_107}; // @[offreg.scala 59:15:@22.4]
  assign _T_113 = $signed(_T_99) + $signed(_GEN_0); // @[offreg.scala 59:15:@22.4]
  assign _T_114 = $signed(_T_99) + $signed(_GEN_0); // @[offreg.scala 59:15:@23.4]
  assign _T_115 = $signed(_T_114); // @[offreg.scala 59:15:@24.4]
  assign _GEN_1 = {{9{_T_112[22]}},_T_112}; // @[offreg.scala 60:15:@25.4]
  assign _T_116 = $signed(_T_100) + $signed(_GEN_1); // @[offreg.scala 60:15:@25.4]
  assign _T_117 = $signed(_T_100) + $signed(_GEN_1); // @[offreg.scala 60:15:@26.4]
  assign _T_118 = $signed(_T_117); // @[offreg.scala 60:15:@27.4]
  assign _T_121 = $signed(_T_104) * $signed(28'sh1); // @[offreg.scala 65:32:@30.4]
  assign _T_122 = $signed(_T_121); // @[offreg.scala 65:52:@31.4]
  assign _T_123 = _T_122[29:6]; // @[offreg.scala 65:60:@32.4]
  assign _T_126 = $signed(_T_109) * $signed(28'sh1); // @[offreg.scala 66:32:@35.4]
  assign _T_127 = $signed(_T_126); // @[offreg.scala 66:52:@36.4]
  assign _T_128 = _T_127[29:6]; // @[offreg.scala 66:60:@37.4]
  assign _GEN_2 = {{8{_T_123[23]}},_T_123}; // @[offreg.scala 59:15:@38.4]
  assign _T_129 = $signed(_T_99) + $signed(_GEN_2); // @[offreg.scala 59:15:@38.4]
  assign _T_130 = $signed(_T_99) + $signed(_GEN_2); // @[offreg.scala 59:15:@39.4]
  assign _T_131 = $signed(_T_130); // @[offreg.scala 59:15:@40.4]
  assign _GEN_3 = {{8{_T_128[23]}},_T_128}; // @[offreg.scala 60:15:@41.4]
  assign _T_132 = $signed(_T_100) + $signed(_GEN_3); // @[offreg.scala 60:15:@41.4]
  assign _T_133 = $signed(_T_100) + $signed(_GEN_3); // @[offreg.scala 60:15:@42.4]
  assign _T_134 = $signed(_T_133); // @[offreg.scala 60:15:@43.4]
  assign _T_137 = $signed(_T_104) * $signed(28'sh2); // @[offreg.scala 65:32:@46.4]
  assign _T_138 = $signed(_T_137); // @[offreg.scala 65:52:@47.4]
  assign _T_139 = _T_138[30:6]; // @[offreg.scala 65:60:@48.4]
  assign _T_142 = $signed(_T_109) * $signed(28'sh2); // @[offreg.scala 66:32:@51.4]
  assign _T_143 = $signed(_T_142); // @[offreg.scala 66:52:@52.4]
  assign _T_144 = _T_143[30:6]; // @[offreg.scala 66:60:@53.4]
  assign _GEN_4 = {{7{_T_139[24]}},_T_139}; // @[offreg.scala 59:15:@54.4]
  assign _T_145 = $signed(_T_99) + $signed(_GEN_4); // @[offreg.scala 59:15:@54.4]
  assign _T_146 = $signed(_T_99) + $signed(_GEN_4); // @[offreg.scala 59:15:@55.4]
  assign _T_147 = $signed(_T_146); // @[offreg.scala 59:15:@56.4]
  assign _GEN_5 = {{7{_T_144[24]}},_T_144}; // @[offreg.scala 60:15:@57.4]
  assign _T_148 = $signed(_T_100) + $signed(_GEN_5); // @[offreg.scala 60:15:@57.4]
  assign _T_149 = $signed(_T_100) + $signed(_GEN_5); // @[offreg.scala 60:15:@58.4]
  assign _T_150 = $signed(_T_149); // @[offreg.scala 60:15:@59.4]
  assign _T_153 = $signed(_T_104) * $signed(28'sh3); // @[offreg.scala 65:32:@62.4]
  assign _T_154 = $signed(_T_153); // @[offreg.scala 65:52:@63.4]
  assign _T_155 = _T_154[30:6]; // @[offreg.scala 65:60:@64.4]
  assign _T_158 = $signed(_T_109) * $signed(28'sh3); // @[offreg.scala 66:32:@67.4]
  assign _T_159 = $signed(_T_158); // @[offreg.scala 66:52:@68.4]
  assign _T_160 = _T_159[30:6]; // @[offreg.scala 66:60:@69.4]
  assign _GEN_6 = {{7{_T_155[24]}},_T_155}; // @[offreg.scala 59:15:@70.4]
  assign _T_161 = $signed(_T_99) + $signed(_GEN_6); // @[offreg.scala 59:15:@70.4]
  assign _T_162 = $signed(_T_99) + $signed(_GEN_6); // @[offreg.scala 59:15:@71.4]
  assign _T_163 = $signed(_T_162); // @[offreg.scala 59:15:@72.4]
  assign _GEN_7 = {{7{_T_160[24]}},_T_160}; // @[offreg.scala 60:15:@73.4]
  assign _T_164 = $signed(_T_100) + $signed(_GEN_7); // @[offreg.scala 60:15:@73.4]
  assign _T_165 = $signed(_T_100) + $signed(_GEN_7); // @[offreg.scala 60:15:@74.4]
  assign _T_166 = $signed(_T_165); // @[offreg.scala 60:15:@75.4]
  assign _T_169 = $signed(_T_104) * $signed(28'sh4); // @[offreg.scala 65:32:@78.4]
  assign _T_170 = $signed(_T_169); // @[offreg.scala 65:52:@79.4]
  assign _T_171 = _T_170[31:6]; // @[offreg.scala 65:60:@80.4]
  assign _T_174 = $signed(_T_109) * $signed(28'sh4); // @[offreg.scala 66:32:@83.4]
  assign _T_175 = $signed(_T_174); // @[offreg.scala 66:52:@84.4]
  assign _T_176 = _T_175[31:6]; // @[offreg.scala 66:60:@85.4]
  assign _GEN_8 = {{6{_T_171[25]}},_T_171}; // @[offreg.scala 59:15:@86.4]
  assign _T_177 = $signed(_T_99) + $signed(_GEN_8); // @[offreg.scala 59:15:@86.4]
  assign _T_178 = $signed(_T_99) + $signed(_GEN_8); // @[offreg.scala 59:15:@87.4]
  assign _T_179 = $signed(_T_178); // @[offreg.scala 59:15:@88.4]
  assign _GEN_9 = {{6{_T_176[25]}},_T_176}; // @[offreg.scala 60:15:@89.4]
  assign _T_180 = $signed(_T_100) + $signed(_GEN_9); // @[offreg.scala 60:15:@89.4]
  assign _T_181 = $signed(_T_100) + $signed(_GEN_9); // @[offreg.scala 60:15:@90.4]
  assign _T_182 = $signed(_T_181); // @[offreg.scala 60:15:@91.4]
  assign _T_185 = $signed(_T_104) * $signed(28'sh5); // @[offreg.scala 65:32:@94.4]
  assign _T_186 = $signed(_T_185); // @[offreg.scala 65:52:@95.4]
  assign _T_187 = _T_186[31:6]; // @[offreg.scala 65:60:@96.4]
  assign _T_190 = $signed(_T_109) * $signed(28'sh5); // @[offreg.scala 66:32:@99.4]
  assign _T_191 = $signed(_T_190); // @[offreg.scala 66:52:@100.4]
  assign _T_192 = _T_191[31:6]; // @[offreg.scala 66:60:@101.4]
  assign _GEN_10 = {{6{_T_187[25]}},_T_187}; // @[offreg.scala 59:15:@102.4]
  assign _T_193 = $signed(_T_99) + $signed(_GEN_10); // @[offreg.scala 59:15:@102.4]
  assign _T_194 = $signed(_T_99) + $signed(_GEN_10); // @[offreg.scala 59:15:@103.4]
  assign _T_195 = $signed(_T_194); // @[offreg.scala 59:15:@104.4]
  assign _GEN_11 = {{6{_T_192[25]}},_T_192}; // @[offreg.scala 60:15:@105.4]
  assign _T_196 = $signed(_T_100) + $signed(_GEN_11); // @[offreg.scala 60:15:@105.4]
  assign _T_197 = $signed(_T_100) + $signed(_GEN_11); // @[offreg.scala 60:15:@106.4]
  assign _T_198 = $signed(_T_197); // @[offreg.scala 60:15:@107.4]
  assign _T_201 = $signed(_T_104) * $signed(28'sh6); // @[offreg.scala 65:32:@110.4]
  assign _T_202 = $signed(_T_201); // @[offreg.scala 65:52:@111.4]
  assign _T_203 = _T_202[31:6]; // @[offreg.scala 65:60:@112.4]
  assign _T_206 = $signed(_T_109) * $signed(28'sh6); // @[offreg.scala 66:32:@115.4]
  assign _T_207 = $signed(_T_206); // @[offreg.scala 66:52:@116.4]
  assign _T_208 = _T_207[31:6]; // @[offreg.scala 66:60:@117.4]
  assign _GEN_12 = {{6{_T_203[25]}},_T_203}; // @[offreg.scala 59:15:@118.4]
  assign _T_209 = $signed(_T_99) + $signed(_GEN_12); // @[offreg.scala 59:15:@118.4]
  assign _T_210 = $signed(_T_99) + $signed(_GEN_12); // @[offreg.scala 59:15:@119.4]
  assign _T_211 = $signed(_T_210); // @[offreg.scala 59:15:@120.4]
  assign _GEN_13 = {{6{_T_208[25]}},_T_208}; // @[offreg.scala 60:15:@121.4]
  assign _T_212 = $signed(_T_100) + $signed(_GEN_13); // @[offreg.scala 60:15:@121.4]
  assign _T_213 = $signed(_T_100) + $signed(_GEN_13); // @[offreg.scala 60:15:@122.4]
  assign _T_214 = $signed(_T_213); // @[offreg.scala 60:15:@123.4]
  assign _T_217 = $signed(_T_104) * $signed(28'sh7); // @[offreg.scala 65:32:@126.4]
  assign _T_218 = $signed(_T_217); // @[offreg.scala 65:52:@127.4]
  assign _T_219 = _T_218[31:6]; // @[offreg.scala 65:60:@128.4]
  assign _T_222 = $signed(_T_109) * $signed(28'sh7); // @[offreg.scala 66:32:@131.4]
  assign _T_223 = $signed(_T_222); // @[offreg.scala 66:52:@132.4]
  assign _T_224 = _T_223[31:6]; // @[offreg.scala 66:60:@133.4]
  assign _GEN_14 = {{6{_T_219[25]}},_T_219}; // @[offreg.scala 59:15:@134.4]
  assign _T_225 = $signed(_T_99) + $signed(_GEN_14); // @[offreg.scala 59:15:@134.4]
  assign _T_226 = $signed(_T_99) + $signed(_GEN_14); // @[offreg.scala 59:15:@135.4]
  assign _T_227 = $signed(_T_226); // @[offreg.scala 59:15:@136.4]
  assign _GEN_15 = {{6{_T_224[25]}},_T_224}; // @[offreg.scala 60:15:@137.4]
  assign _T_228 = $signed(_T_100) + $signed(_GEN_15); // @[offreg.scala 60:15:@137.4]
  assign _T_229 = $signed(_T_100) + $signed(_GEN_15); // @[offreg.scala 60:15:@138.4]
  assign _T_230 = $signed(_T_229); // @[offreg.scala 60:15:@139.4]
  assign _T_233 = $signed(_T_104) * $signed(28'sh8); // @[offreg.scala 65:32:@142.4]
  assign _T_234 = $signed(_T_233); // @[offreg.scala 65:52:@143.4]
  assign _T_235 = _T_234[32:6]; // @[offreg.scala 65:60:@144.4]
  assign _T_238 = $signed(_T_109) * $signed(28'sh8); // @[offreg.scala 66:32:@147.4]
  assign _T_239 = $signed(_T_238); // @[offreg.scala 66:52:@148.4]
  assign _T_240 = _T_239[32:6]; // @[offreg.scala 66:60:@149.4]
  assign _GEN_16 = {{5{_T_235[26]}},_T_235}; // @[offreg.scala 59:15:@150.4]
  assign _T_241 = $signed(_T_99) + $signed(_GEN_16); // @[offreg.scala 59:15:@150.4]
  assign _T_242 = $signed(_T_99) + $signed(_GEN_16); // @[offreg.scala 59:15:@151.4]
  assign _T_243 = $signed(_T_242); // @[offreg.scala 59:15:@152.4]
  assign _GEN_17 = {{5{_T_240[26]}},_T_240}; // @[offreg.scala 60:15:@153.4]
  assign _T_244 = $signed(_T_100) + $signed(_GEN_17); // @[offreg.scala 60:15:@153.4]
  assign _T_245 = $signed(_T_100) + $signed(_GEN_17); // @[offreg.scala 60:15:@154.4]
  assign _T_246 = $signed(_T_245); // @[offreg.scala 60:15:@155.4]
  assign _T_249 = $signed(_T_104) * $signed(28'sh9); // @[offreg.scala 65:32:@158.4]
  assign _T_250 = $signed(_T_249); // @[offreg.scala 65:52:@159.4]
  assign _T_251 = _T_250[32:6]; // @[offreg.scala 65:60:@160.4]
  assign _T_254 = $signed(_T_109) * $signed(28'sh9); // @[offreg.scala 66:32:@163.4]
  assign _T_255 = $signed(_T_254); // @[offreg.scala 66:52:@164.4]
  assign _T_256 = _T_255[32:6]; // @[offreg.scala 66:60:@165.4]
  assign _GEN_18 = {{5{_T_251[26]}},_T_251}; // @[offreg.scala 59:15:@166.4]
  assign _T_257 = $signed(_T_99) + $signed(_GEN_18); // @[offreg.scala 59:15:@166.4]
  assign _T_258 = $signed(_T_99) + $signed(_GEN_18); // @[offreg.scala 59:15:@167.4]
  assign _T_259 = $signed(_T_258); // @[offreg.scala 59:15:@168.4]
  assign _GEN_19 = {{5{_T_256[26]}},_T_256}; // @[offreg.scala 60:15:@169.4]
  assign _T_260 = $signed(_T_100) + $signed(_GEN_19); // @[offreg.scala 60:15:@169.4]
  assign _T_261 = $signed(_T_100) + $signed(_GEN_19); // @[offreg.scala 60:15:@170.4]
  assign _T_262 = $signed(_T_261); // @[offreg.scala 60:15:@171.4]
  assign _T_265 = $signed(_T_104) * $signed(28'sha); // @[offreg.scala 65:32:@174.4]
  assign _T_266 = $signed(_T_265); // @[offreg.scala 65:52:@175.4]
  assign _T_267 = _T_266[32:6]; // @[offreg.scala 65:60:@176.4]
  assign _T_270 = $signed(_T_109) * $signed(28'sha); // @[offreg.scala 66:32:@179.4]
  assign _T_271 = $signed(_T_270); // @[offreg.scala 66:52:@180.4]
  assign _T_272 = _T_271[32:6]; // @[offreg.scala 66:60:@181.4]
  assign _GEN_20 = {{5{_T_267[26]}},_T_267}; // @[offreg.scala 59:15:@182.4]
  assign _T_273 = $signed(_T_99) + $signed(_GEN_20); // @[offreg.scala 59:15:@182.4]
  assign _T_274 = $signed(_T_99) + $signed(_GEN_20); // @[offreg.scala 59:15:@183.4]
  assign _T_275 = $signed(_T_274); // @[offreg.scala 59:15:@184.4]
  assign _GEN_21 = {{5{_T_272[26]}},_T_272}; // @[offreg.scala 60:15:@185.4]
  assign _T_276 = $signed(_T_100) + $signed(_GEN_21); // @[offreg.scala 60:15:@185.4]
  assign _T_277 = $signed(_T_100) + $signed(_GEN_21); // @[offreg.scala 60:15:@186.4]
  assign _T_278 = $signed(_T_277); // @[offreg.scala 60:15:@187.4]
  assign _T_281 = $signed(_T_104) * $signed(28'shb); // @[offreg.scala 65:32:@190.4]
  assign _T_282 = $signed(_T_281); // @[offreg.scala 65:52:@191.4]
  assign _T_283 = _T_282[32:6]; // @[offreg.scala 65:60:@192.4]
  assign _T_286 = $signed(_T_109) * $signed(28'shb); // @[offreg.scala 66:32:@195.4]
  assign _T_287 = $signed(_T_286); // @[offreg.scala 66:52:@196.4]
  assign _T_288 = _T_287[32:6]; // @[offreg.scala 66:60:@197.4]
  assign _GEN_22 = {{5{_T_283[26]}},_T_283}; // @[offreg.scala 59:15:@198.4]
  assign _T_289 = $signed(_T_99) + $signed(_GEN_22); // @[offreg.scala 59:15:@198.4]
  assign _T_290 = $signed(_T_99) + $signed(_GEN_22); // @[offreg.scala 59:15:@199.4]
  assign _T_291 = $signed(_T_290); // @[offreg.scala 59:15:@200.4]
  assign _GEN_23 = {{5{_T_288[26]}},_T_288}; // @[offreg.scala 60:15:@201.4]
  assign _T_292 = $signed(_T_100) + $signed(_GEN_23); // @[offreg.scala 60:15:@201.4]
  assign _T_293 = $signed(_T_100) + $signed(_GEN_23); // @[offreg.scala 60:15:@202.4]
  assign _T_294 = $signed(_T_293); // @[offreg.scala 60:15:@203.4]
  assign _T_297 = $signed(_T_104) * $signed(28'shc); // @[offreg.scala 65:32:@206.4]
  assign _T_298 = $signed(_T_297); // @[offreg.scala 65:52:@207.4]
  assign _T_299 = _T_298[32:6]; // @[offreg.scala 65:60:@208.4]
  assign _T_302 = $signed(_T_109) * $signed(28'shc); // @[offreg.scala 66:32:@211.4]
  assign _T_303 = $signed(_T_302); // @[offreg.scala 66:52:@212.4]
  assign _T_304 = _T_303[32:6]; // @[offreg.scala 66:60:@213.4]
  assign _GEN_24 = {{5{_T_299[26]}},_T_299}; // @[offreg.scala 59:15:@214.4]
  assign _T_305 = $signed(_T_99) + $signed(_GEN_24); // @[offreg.scala 59:15:@214.4]
  assign _T_306 = $signed(_T_99) + $signed(_GEN_24); // @[offreg.scala 59:15:@215.4]
  assign _T_307 = $signed(_T_306); // @[offreg.scala 59:15:@216.4]
  assign _GEN_25 = {{5{_T_304[26]}},_T_304}; // @[offreg.scala 60:15:@217.4]
  assign _T_308 = $signed(_T_100) + $signed(_GEN_25); // @[offreg.scala 60:15:@217.4]
  assign _T_309 = $signed(_T_100) + $signed(_GEN_25); // @[offreg.scala 60:15:@218.4]
  assign _T_310 = $signed(_T_309); // @[offreg.scala 60:15:@219.4]
  assign _T_313 = $signed(_T_104) * $signed(28'shd); // @[offreg.scala 65:32:@222.4]
  assign _T_314 = $signed(_T_313); // @[offreg.scala 65:52:@223.4]
  assign _T_315 = _T_314[32:6]; // @[offreg.scala 65:60:@224.4]
  assign _T_318 = $signed(_T_109) * $signed(28'shd); // @[offreg.scala 66:32:@227.4]
  assign _T_319 = $signed(_T_318); // @[offreg.scala 66:52:@228.4]
  assign _T_320 = _T_319[32:6]; // @[offreg.scala 66:60:@229.4]
  assign _GEN_26 = {{5{_T_315[26]}},_T_315}; // @[offreg.scala 59:15:@230.4]
  assign _T_321 = $signed(_T_99) + $signed(_GEN_26); // @[offreg.scala 59:15:@230.4]
  assign _T_322 = $signed(_T_99) + $signed(_GEN_26); // @[offreg.scala 59:15:@231.4]
  assign _T_323 = $signed(_T_322); // @[offreg.scala 59:15:@232.4]
  assign _GEN_27 = {{5{_T_320[26]}},_T_320}; // @[offreg.scala 60:15:@233.4]
  assign _T_324 = $signed(_T_100) + $signed(_GEN_27); // @[offreg.scala 60:15:@233.4]
  assign _T_325 = $signed(_T_100) + $signed(_GEN_27); // @[offreg.scala 60:15:@234.4]
  assign _T_326 = $signed(_T_325); // @[offreg.scala 60:15:@235.4]
  assign _T_329 = $signed(_T_104) * $signed(28'she); // @[offreg.scala 65:32:@238.4]
  assign _T_330 = $signed(_T_329); // @[offreg.scala 65:52:@239.4]
  assign _T_331 = _T_330[32:6]; // @[offreg.scala 65:60:@240.4]
  assign _T_334 = $signed(_T_109) * $signed(28'she); // @[offreg.scala 66:32:@243.4]
  assign _T_335 = $signed(_T_334); // @[offreg.scala 66:52:@244.4]
  assign _T_336 = _T_335[32:6]; // @[offreg.scala 66:60:@245.4]
  assign _GEN_28 = {{5{_T_331[26]}},_T_331}; // @[offreg.scala 59:15:@246.4]
  assign _T_337 = $signed(_T_99) + $signed(_GEN_28); // @[offreg.scala 59:15:@246.4]
  assign _T_338 = $signed(_T_99) + $signed(_GEN_28); // @[offreg.scala 59:15:@247.4]
  assign _T_339 = $signed(_T_338); // @[offreg.scala 59:15:@248.4]
  assign _GEN_29 = {{5{_T_336[26]}},_T_336}; // @[offreg.scala 60:15:@249.4]
  assign _T_340 = $signed(_T_100) + $signed(_GEN_29); // @[offreg.scala 60:15:@249.4]
  assign _T_341 = $signed(_T_100) + $signed(_GEN_29); // @[offreg.scala 60:15:@250.4]
  assign _T_342 = $signed(_T_341); // @[offreg.scala 60:15:@251.4]
  assign _T_345 = $signed(_T_104) * $signed(28'shf); // @[offreg.scala 65:32:@254.4]
  assign _T_346 = $signed(_T_345); // @[offreg.scala 65:52:@255.4]
  assign _T_347 = _T_346[32:6]; // @[offreg.scala 65:60:@256.4]
  assign _T_350 = $signed(_T_109) * $signed(28'shf); // @[offreg.scala 66:32:@259.4]
  assign _T_351 = $signed(_T_350); // @[offreg.scala 66:52:@260.4]
  assign _T_352 = _T_351[32:6]; // @[offreg.scala 66:60:@261.4]
  assign _GEN_30 = {{5{_T_347[26]}},_T_347}; // @[offreg.scala 59:15:@262.4]
  assign _T_353 = $signed(_T_99) + $signed(_GEN_30); // @[offreg.scala 59:15:@262.4]
  assign _T_354 = $signed(_T_99) + $signed(_GEN_30); // @[offreg.scala 59:15:@263.4]
  assign _T_355 = $signed(_T_354); // @[offreg.scala 59:15:@264.4]
  assign _GEN_31 = {{5{_T_352[26]}},_T_352}; // @[offreg.scala 60:15:@265.4]
  assign _T_356 = $signed(_T_100) + $signed(_GEN_31); // @[offreg.scala 60:15:@265.4]
  assign _T_357 = $signed(_T_100) + $signed(_GEN_31); // @[offreg.scala 60:15:@266.4]
  assign _T_358 = $signed(_T_357); // @[offreg.scala 60:15:@267.4]
  assign _T_393 = $signed(_T_99) + $signed(32'sh1000000); // @[offreg.scala 59:15:@332.4]
  assign _T_394 = $signed(_T_99) + $signed(32'sh1000000); // @[offreg.scala 59:15:@333.4]
  assign _T_395 = $signed(_T_394); // @[offreg.scala 59:15:@334.4]
  assign _T_396 = $signed(_T_100) + $signed(32'sh600000); // @[offreg.scala 60:15:@335.4]
  assign _T_397 = $signed(_T_100) + $signed(32'sh600000); // @[offreg.scala 60:15:@336.4]
  assign _T_398 = $signed(_T_397); // @[offreg.scala 60:15:@337.4]
  assign _T_399 = $signed(_T_115) < $signed(_T_395); // @[offreg.scala 70:12:@338.4]
  assign _T_400 = $signed(_T_118) < $signed(_T_398); // @[offreg.scala 70:26:@339.4]
  assign vld_0 = _T_399 & _T_400; // @[offreg.scala 70:20:@340.4]
  assign _T_401 = $signed(_T_131) < $signed(_T_395); // @[offreg.scala 70:12:@341.4]
  assign _T_402 = $signed(_T_134) < $signed(_T_398); // @[offreg.scala 70:26:@342.4]
  assign vld_1 = _T_401 & _T_402; // @[offreg.scala 70:20:@343.4]
  assign _T_403 = $signed(_T_147) < $signed(_T_395); // @[offreg.scala 70:12:@344.4]
  assign _T_404 = $signed(_T_150) < $signed(_T_398); // @[offreg.scala 70:26:@345.4]
  assign vld_2 = _T_403 & _T_404; // @[offreg.scala 70:20:@346.4]
  assign _T_405 = $signed(_T_163) < $signed(_T_395); // @[offreg.scala 70:12:@347.4]
  assign _T_406 = $signed(_T_166) < $signed(_T_398); // @[offreg.scala 70:26:@348.4]
  assign vld_3 = _T_405 & _T_406; // @[offreg.scala 70:20:@349.4]
  assign _T_407 = $signed(_T_179) < $signed(_T_395); // @[offreg.scala 70:12:@350.4]
  assign _T_408 = $signed(_T_182) < $signed(_T_398); // @[offreg.scala 70:26:@351.4]
  assign vld_4 = _T_407 & _T_408; // @[offreg.scala 70:20:@352.4]
  assign _T_409 = $signed(_T_195) < $signed(_T_395); // @[offreg.scala 70:12:@353.4]
  assign _T_410 = $signed(_T_198) < $signed(_T_398); // @[offreg.scala 70:26:@354.4]
  assign vld_5 = _T_409 & _T_410; // @[offreg.scala 70:20:@355.4]
  assign _T_411 = $signed(_T_211) < $signed(_T_395); // @[offreg.scala 70:12:@356.4]
  assign _T_412 = $signed(_T_214) < $signed(_T_398); // @[offreg.scala 70:26:@357.4]
  assign vld_6 = _T_411 & _T_412; // @[offreg.scala 70:20:@358.4]
  assign _T_413 = $signed(_T_227) < $signed(_T_395); // @[offreg.scala 70:12:@359.4]
  assign _T_414 = $signed(_T_230) < $signed(_T_398); // @[offreg.scala 70:26:@360.4]
  assign vld_7 = _T_413 & _T_414; // @[offreg.scala 70:20:@361.4]
  assign _T_415 = $signed(_T_243) < $signed(_T_395); // @[offreg.scala 70:12:@362.4]
  assign _T_416 = $signed(_T_246) < $signed(_T_398); // @[offreg.scala 70:26:@363.4]
  assign vld_8 = _T_415 & _T_416; // @[offreg.scala 70:20:@364.4]
  assign _T_417 = $signed(_T_259) < $signed(_T_395); // @[offreg.scala 70:12:@365.4]
  assign _T_418 = $signed(_T_262) < $signed(_T_398); // @[offreg.scala 70:26:@366.4]
  assign vld_9 = _T_417 & _T_418; // @[offreg.scala 70:20:@367.4]
  assign _T_419 = $signed(_T_275) < $signed(_T_395); // @[offreg.scala 70:12:@368.4]
  assign _T_420 = $signed(_T_278) < $signed(_T_398); // @[offreg.scala 70:26:@369.4]
  assign vld_10 = _T_419 & _T_420; // @[offreg.scala 70:20:@370.4]
  assign _T_421 = $signed(_T_291) < $signed(_T_395); // @[offreg.scala 70:12:@371.4]
  assign _T_422 = $signed(_T_294) < $signed(_T_398); // @[offreg.scala 70:26:@372.4]
  assign vld_11 = _T_421 & _T_422; // @[offreg.scala 70:20:@373.4]
  assign _T_423 = $signed(_T_307) < $signed(_T_395); // @[offreg.scala 70:12:@374.4]
  assign _T_424 = $signed(_T_310) < $signed(_T_398); // @[offreg.scala 70:26:@375.4]
  assign vld_12 = _T_423 & _T_424; // @[offreg.scala 70:20:@376.4]
  assign _T_425 = $signed(_T_323) < $signed(_T_395); // @[offreg.scala 70:12:@377.4]
  assign _T_426 = $signed(_T_326) < $signed(_T_398); // @[offreg.scala 70:26:@378.4]
  assign vld_13 = _T_425 & _T_426; // @[offreg.scala 70:20:@379.4]
  assign _T_427 = $signed(_T_339) < $signed(_T_395); // @[offreg.scala 70:12:@380.4]
  assign _T_428 = $signed(_T_342) < $signed(_T_398); // @[offreg.scala 70:26:@381.4]
  assign vld_14 = _T_427 & _T_428; // @[offreg.scala 70:20:@382.4]
  assign _T_429 = $signed(_T_355) < $signed(_T_395); // @[offreg.scala 70:12:@383.4]
  assign _T_430 = $signed(_T_358) < $signed(_T_398); // @[offreg.scala 70:26:@384.4]
  assign vld_15 = _T_429 & _T_430; // @[offreg.scala 70:20:@385.4]
  assign _GEN_32 = {{1'd0}, vld_1}; // @[offreg.scala 32:52:@387.4]
  assign _T_432 = _GEN_32 << 1; // @[offreg.scala 32:52:@387.4]
  assign _GEN_33 = {{2'd0}, vld_2}; // @[offreg.scala 32:52:@388.4]
  assign _T_433 = _GEN_33 << 2; // @[offreg.scala 32:52:@388.4]
  assign _GEN_34 = {{3'd0}, vld_3}; // @[offreg.scala 32:52:@389.4]
  assign _T_434 = _GEN_34 << 3; // @[offreg.scala 32:52:@389.4]
  assign _GEN_35 = {{4'd0}, vld_4}; // @[offreg.scala 32:52:@390.4]
  assign _T_435 = _GEN_35 << 4; // @[offreg.scala 32:52:@390.4]
  assign _GEN_36 = {{5'd0}, vld_5}; // @[offreg.scala 32:52:@391.4]
  assign _T_436 = _GEN_36 << 5; // @[offreg.scala 32:52:@391.4]
  assign _GEN_37 = {{6'd0}, vld_6}; // @[offreg.scala 32:52:@392.4]
  assign _T_437 = _GEN_37 << 6; // @[offreg.scala 32:52:@392.4]
  assign _GEN_38 = {{7'd0}, vld_7}; // @[offreg.scala 32:52:@393.4]
  assign _T_438 = _GEN_38 << 7; // @[offreg.scala 32:52:@393.4]
  assign _GEN_39 = {{8'd0}, vld_8}; // @[offreg.scala 32:52:@394.4]
  assign _T_439 = _GEN_39 << 8; // @[offreg.scala 32:52:@394.4]
  assign _GEN_40 = {{9'd0}, vld_9}; // @[offreg.scala 32:52:@395.4]
  assign _T_440 = _GEN_40 << 9; // @[offreg.scala 32:52:@395.4]
  assign _GEN_41 = {{10'd0}, vld_10}; // @[offreg.scala 32:52:@396.4]
  assign _T_441 = _GEN_41 << 10; // @[offreg.scala 32:52:@396.4]
  assign _GEN_42 = {{11'd0}, vld_11}; // @[offreg.scala 32:52:@397.4]
  assign _T_442 = _GEN_42 << 11; // @[offreg.scala 32:52:@397.4]
  assign _GEN_43 = {{12'd0}, vld_12}; // @[offreg.scala 32:52:@398.4]
  assign _T_443 = _GEN_43 << 12; // @[offreg.scala 32:52:@398.4]
  assign _GEN_44 = {{13'd0}, vld_13}; // @[offreg.scala 32:52:@399.4]
  assign _T_444 = _GEN_44 << 13; // @[offreg.scala 32:52:@399.4]
  assign _GEN_45 = {{14'd0}, vld_14}; // @[offreg.scala 32:52:@400.4]
  assign _T_445 = _GEN_45 << 14; // @[offreg.scala 32:52:@400.4]
  assign _GEN_46 = {{15'd0}, vld_15}; // @[offreg.scala 32:52:@401.4]
  assign _T_446 = _GEN_46 << 15; // @[offreg.scala 32:52:@401.4]
  assign _GEN_47 = {{1'd0}, vld_0}; // @[offreg.scala 32:74:@403.4]
  assign _T_449 = _GEN_47 | _T_432; // @[offreg.scala 32:74:@403.4]
  assign _GEN_48 = {{1'd0}, _T_449}; // @[offreg.scala 32:74:@404.4]
  assign _T_450 = _GEN_48 | _T_433; // @[offreg.scala 32:74:@404.4]
  assign _GEN_49 = {{1'd0}, _T_450}; // @[offreg.scala 32:74:@405.4]
  assign _T_451 = _GEN_49 | _T_434; // @[offreg.scala 32:74:@405.4]
  assign _GEN_50 = {{1'd0}, _T_451}; // @[offreg.scala 32:74:@406.4]
  assign _T_452 = _GEN_50 | _T_435; // @[offreg.scala 32:74:@406.4]
  assign _GEN_51 = {{1'd0}, _T_452}; // @[offreg.scala 32:74:@407.4]
  assign _T_453 = _GEN_51 | _T_436; // @[offreg.scala 32:74:@407.4]
  assign _GEN_52 = {{1'd0}, _T_453}; // @[offreg.scala 32:74:@408.4]
  assign _T_454 = _GEN_52 | _T_437; // @[offreg.scala 32:74:@408.4]
  assign _GEN_53 = {{1'd0}, _T_454}; // @[offreg.scala 32:74:@409.4]
  assign _T_455 = _GEN_53 | _T_438; // @[offreg.scala 32:74:@409.4]
  assign _GEN_54 = {{1'd0}, _T_455}; // @[offreg.scala 32:74:@410.4]
  assign _T_456 = _GEN_54 | _T_439; // @[offreg.scala 32:74:@410.4]
  assign _GEN_55 = {{1'd0}, _T_456}; // @[offreg.scala 32:74:@411.4]
  assign _T_457 = _GEN_55 | _T_440; // @[offreg.scala 32:74:@411.4]
  assign _GEN_56 = {{1'd0}, _T_457}; // @[offreg.scala 32:74:@412.4]
  assign _T_458 = _GEN_56 | _T_441; // @[offreg.scala 32:74:@412.4]
  assign _GEN_57 = {{1'd0}, _T_458}; // @[offreg.scala 32:74:@413.4]
  assign _T_459 = _GEN_57 | _T_442; // @[offreg.scala 32:74:@413.4]
  assign _GEN_58 = {{1'd0}, _T_459}; // @[offreg.scala 32:74:@414.4]
  assign _T_460 = _GEN_58 | _T_443; // @[offreg.scala 32:74:@414.4]
  assign _GEN_59 = {{1'd0}, _T_460}; // @[offreg.scala 32:74:@415.4]
  assign _T_461 = _GEN_59 | _T_444; // @[offreg.scala 32:74:@415.4]
  assign _GEN_60 = {{1'd0}, _T_461}; // @[offreg.scala 32:74:@416.4]
  assign _T_462 = _GEN_60 | _T_445; // @[offreg.scala 32:74:@416.4]
  assign _GEN_61 = {{1'd0}, _T_462}; // @[offreg.scala 32:74:@417.4]
  assign _T_463 = _GEN_61 | _T_446; // @[offreg.scala 32:74:@417.4]
  assign io_offset_x_0 = $signed(_T_115); // @[offreg.scala 27:17:@284.4]
  assign io_offset_x_1 = $signed(_T_131); // @[offreg.scala 27:17:@285.4]
  assign io_offset_x_2 = $signed(_T_147); // @[offreg.scala 27:17:@286.4]
  assign io_offset_x_3 = $signed(_T_163); // @[offreg.scala 27:17:@287.4]
  assign io_offset_x_4 = $signed(_T_179); // @[offreg.scala 27:17:@288.4]
  assign io_offset_x_5 = $signed(_T_195); // @[offreg.scala 27:17:@289.4]
  assign io_offset_x_6 = $signed(_T_211); // @[offreg.scala 27:17:@290.4]
  assign io_offset_x_7 = $signed(_T_227); // @[offreg.scala 27:17:@291.4]
  assign io_offset_x_8 = $signed(_T_243); // @[offreg.scala 27:17:@292.4]
  assign io_offset_x_9 = $signed(_T_259); // @[offreg.scala 27:17:@293.4]
  assign io_offset_x_10 = $signed(_T_275); // @[offreg.scala 27:17:@294.4]
  assign io_offset_x_11 = $signed(_T_291); // @[offreg.scala 27:17:@295.4]
  assign io_offset_x_12 = $signed(_T_307); // @[offreg.scala 27:17:@296.4]
  assign io_offset_x_13 = $signed(_T_323); // @[offreg.scala 27:17:@297.4]
  assign io_offset_x_14 = $signed(_T_339); // @[offreg.scala 27:17:@298.4]
  assign io_offset_x_15 = $signed(_T_355); // @[offreg.scala 27:17:@299.4]
  assign io_offset_y_0 = $signed(_T_118); // @[offreg.scala 28:17:@316.4]
  assign io_offset_y_1 = $signed(_T_134); // @[offreg.scala 28:17:@317.4]
  assign io_offset_y_2 = $signed(_T_150); // @[offreg.scala 28:17:@318.4]
  assign io_offset_y_3 = $signed(_T_166); // @[offreg.scala 28:17:@319.4]
  assign io_offset_y_4 = $signed(_T_182); // @[offreg.scala 28:17:@320.4]
  assign io_offset_y_5 = $signed(_T_198); // @[offreg.scala 28:17:@321.4]
  assign io_offset_y_6 = $signed(_T_214); // @[offreg.scala 28:17:@322.4]
  assign io_offset_y_7 = $signed(_T_230); // @[offreg.scala 28:17:@323.4]
  assign io_offset_y_8 = $signed(_T_246); // @[offreg.scala 28:17:@324.4]
  assign io_offset_y_9 = $signed(_T_262); // @[offreg.scala 28:17:@325.4]
  assign io_offset_y_10 = $signed(_T_278); // @[offreg.scala 28:17:@326.4]
  assign io_offset_y_11 = $signed(_T_294); // @[offreg.scala 28:17:@327.4]
  assign io_offset_y_12 = $signed(_T_310); // @[offreg.scala 28:17:@328.4]
  assign io_offset_y_13 = $signed(_T_326); // @[offreg.scala 28:17:@329.4]
  assign io_offset_y_14 = $signed(_T_342); // @[offreg.scala 28:17:@330.4]
  assign io_offset_y_15 = $signed(_T_358); // @[offreg.scala 28:17:@331.4]
  assign io_vld = {{16'd0}, _T_463}; // @[offreg.scala 32:12:@418.4]
endmodule
